
      <head>
        <meta charset="UTF-8">
        <link rel="icon" href="https://fav.farm/💩" />
      </head>
      <p>You should end your url with .svg, like <a href="/cat.svg">/cat.svg</a></p>
      <style>
        body {
          text-align: center;
          font-family: sans-serif;
          height: 100vh;
          display: grid;
          place-items: center;
          font-size: 2em;
        }
      </style>

        